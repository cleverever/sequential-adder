module sequential_adder_tb;
endmodule